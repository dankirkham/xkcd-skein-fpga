module hash_bits_off (
  input [1023:0] hash_xor_i,
  output reg [9:0] bits_off_o
);

always @(*) begin
  bits_off_o = hash_xor_i[0] + hash_xor_i[1] + hash_xor_i[2] + hash_xor_i[3] + hash_xor_i[4] + hash_xor_i[5] + hash_xor_i[6] + hash_xor_i[7] + hash_xor_i[8] + hash_xor_i[9] + hash_xor_i[10] + hash_xor_i[11] + hash_xor_i[12] + hash_xor_i[13] + hash_xor_i[14] + hash_xor_i[15] + hash_xor_i[16] + hash_xor_i[17] + hash_xor_i[18] + hash_xor_i[19] + hash_xor_i[20] + hash_xor_i[21] + hash_xor_i[22] + hash_xor_i[23] + hash_xor_i[24] + hash_xor_i[25] + hash_xor_i[26] + hash_xor_i[27] + hash_xor_i[28] + hash_xor_i[29] + hash_xor_i[30] + hash_xor_i[31] + hash_xor_i[32] + hash_xor_i[33] + hash_xor_i[34] + hash_xor_i[35] + hash_xor_i[36] + hash_xor_i[37] + hash_xor_i[38] + hash_xor_i[39] + hash_xor_i[40] + hash_xor_i[41] + hash_xor_i[42] + hash_xor_i[43] + hash_xor_i[44] + hash_xor_i[45] + hash_xor_i[46] + hash_xor_i[47] + hash_xor_i[48] + hash_xor_i[49] + hash_xor_i[50] + hash_xor_i[51] + hash_xor_i[52] + hash_xor_i[53] + hash_xor_i[54] + hash_xor_i[55] + hash_xor_i[56] + hash_xor_i[57] + hash_xor_i[58] + hash_xor_i[59] + hash_xor_i[60] + hash_xor_i[61] + hash_xor_i[62] + hash_xor_i[63] + hash_xor_i[64] + hash_xor_i[65] + hash_xor_i[66] + hash_xor_i[67] + hash_xor_i[68] + hash_xor_i[69] + hash_xor_i[70] + hash_xor_i[71] + hash_xor_i[72] + hash_xor_i[73] + hash_xor_i[74] + hash_xor_i[75] + hash_xor_i[76] + hash_xor_i[77] + hash_xor_i[78] + hash_xor_i[79] + hash_xor_i[80] + hash_xor_i[81] + hash_xor_i[82] + hash_xor_i[83] + hash_xor_i[84] + hash_xor_i[85] + hash_xor_i[86] + hash_xor_i[87] + hash_xor_i[88] + hash_xor_i[89] + hash_xor_i[90] + hash_xor_i[91] + hash_xor_i[92] + hash_xor_i[93] + hash_xor_i[94] + hash_xor_i[95] + hash_xor_i[96] + hash_xor_i[97] + hash_xor_i[98] + hash_xor_i[99] + hash_xor_i[100] + hash_xor_i[101] + hash_xor_i[102] + hash_xor_i[103] + hash_xor_i[104] + hash_xor_i[105] + hash_xor_i[106] + hash_xor_i[107] + hash_xor_i[108] + hash_xor_i[109] + hash_xor_i[110] + hash_xor_i[111] + hash_xor_i[112] + hash_xor_i[113] + hash_xor_i[114] + hash_xor_i[115] + hash_xor_i[116] + hash_xor_i[117] + hash_xor_i[118] + hash_xor_i[119] + hash_xor_i[120] + hash_xor_i[121] + hash_xor_i[122] + hash_xor_i[123] + hash_xor_i[124] + hash_xor_i[125] + hash_xor_i[126] + hash_xor_i[127] + hash_xor_i[128] + hash_xor_i[129] + hash_xor_i[130] + hash_xor_i[131] + hash_xor_i[132] + hash_xor_i[133] + hash_xor_i[134] + hash_xor_i[135] + hash_xor_i[136] + hash_xor_i[137] + hash_xor_i[138] + hash_xor_i[139] + hash_xor_i[140] + hash_xor_i[141] + hash_xor_i[142] + hash_xor_i[143] + hash_xor_i[144] + hash_xor_i[145] + hash_xor_i[146] + hash_xor_i[147] + hash_xor_i[148] + hash_xor_i[149] + hash_xor_i[150] + hash_xor_i[151] + hash_xor_i[152] + hash_xor_i[153] + hash_xor_i[154] + hash_xor_i[155] + hash_xor_i[156] + hash_xor_i[157] + hash_xor_i[158] + hash_xor_i[159] + hash_xor_i[160] + hash_xor_i[161] + hash_xor_i[162] + hash_xor_i[163] + hash_xor_i[164] + hash_xor_i[165] + hash_xor_i[166] + hash_xor_i[167] + hash_xor_i[168] + hash_xor_i[169] + hash_xor_i[170] + hash_xor_i[171] + hash_xor_i[172] + hash_xor_i[173] + hash_xor_i[174] + hash_xor_i[175] + hash_xor_i[176] + hash_xor_i[177] + hash_xor_i[178] + hash_xor_i[179] + hash_xor_i[180] + hash_xor_i[181] + hash_xor_i[182] + hash_xor_i[183] + hash_xor_i[184] + hash_xor_i[185] + hash_xor_i[186] + hash_xor_i[187] + hash_xor_i[188] + hash_xor_i[189] + hash_xor_i[190] + hash_xor_i[191] + hash_xor_i[192] + hash_xor_i[193] + hash_xor_i[194] + hash_xor_i[195] + hash_xor_i[196] + hash_xor_i[197] + hash_xor_i[198] + hash_xor_i[199] + hash_xor_i[200] + hash_xor_i[201] + hash_xor_i[202] + hash_xor_i[203] + hash_xor_i[204] + hash_xor_i[205] + hash_xor_i[206] + hash_xor_i[207] + hash_xor_i[208] + hash_xor_i[209] + hash_xor_i[210] + hash_xor_i[211] + hash_xor_i[212] + hash_xor_i[213] + hash_xor_i[214] + hash_xor_i[215] + hash_xor_i[216] + hash_xor_i[217] + hash_xor_i[218] + hash_xor_i[219] + hash_xor_i[220] + hash_xor_i[221] + hash_xor_i[222] + hash_xor_i[223] + hash_xor_i[224] + hash_xor_i[225] + hash_xor_i[226] + hash_xor_i[227] + hash_xor_i[228] + hash_xor_i[229] + hash_xor_i[230] + hash_xor_i[231] + hash_xor_i[232] + hash_xor_i[233] + hash_xor_i[234] + hash_xor_i[235] + hash_xor_i[236] + hash_xor_i[237] + hash_xor_i[238] + hash_xor_i[239] + hash_xor_i[240] + hash_xor_i[241] + hash_xor_i[242] + hash_xor_i[243] + hash_xor_i[244] + hash_xor_i[245] + hash_xor_i[246] + hash_xor_i[247] + hash_xor_i[248] + hash_xor_i[249] + hash_xor_i[250] + hash_xor_i[251] + hash_xor_i[252] + hash_xor_i[253] + hash_xor_i[254] + hash_xor_i[255] + hash_xor_i[256] + hash_xor_i[257] + hash_xor_i[258] + hash_xor_i[259] + hash_xor_i[260] + hash_xor_i[261] + hash_xor_i[262] + hash_xor_i[263] + hash_xor_i[264] + hash_xor_i[265] + hash_xor_i[266] + hash_xor_i[267] + hash_xor_i[268] + hash_xor_i[269] + hash_xor_i[270] + hash_xor_i[271] + hash_xor_i[272] + hash_xor_i[273] + hash_xor_i[274] + hash_xor_i[275] + hash_xor_i[276] + hash_xor_i[277] + hash_xor_i[278] + hash_xor_i[279] + hash_xor_i[280] + hash_xor_i[281] + hash_xor_i[282] + hash_xor_i[283] + hash_xor_i[284] + hash_xor_i[285] + hash_xor_i[286] + hash_xor_i[287] + hash_xor_i[288] + hash_xor_i[289] + hash_xor_i[290] + hash_xor_i[291] + hash_xor_i[292] + hash_xor_i[293] + hash_xor_i[294] + hash_xor_i[295] + hash_xor_i[296] + hash_xor_i[297] + hash_xor_i[298] + hash_xor_i[299] + hash_xor_i[300] + hash_xor_i[301] + hash_xor_i[302] + hash_xor_i[303] + hash_xor_i[304] + hash_xor_i[305] + hash_xor_i[306] + hash_xor_i[307] + hash_xor_i[308] + hash_xor_i[309] + hash_xor_i[310] + hash_xor_i[311] + hash_xor_i[312] + hash_xor_i[313] + hash_xor_i[314] + hash_xor_i[315] + hash_xor_i[316] + hash_xor_i[317] + hash_xor_i[318] + hash_xor_i[319] + hash_xor_i[320] + hash_xor_i[321] + hash_xor_i[322] + hash_xor_i[323] + hash_xor_i[324] + hash_xor_i[325] + hash_xor_i[326] + hash_xor_i[327] + hash_xor_i[328] + hash_xor_i[329] + hash_xor_i[330] + hash_xor_i[331] + hash_xor_i[332] + hash_xor_i[333] + hash_xor_i[334] + hash_xor_i[335] + hash_xor_i[336] + hash_xor_i[337] + hash_xor_i[338] + hash_xor_i[339] + hash_xor_i[340] + hash_xor_i[341] + hash_xor_i[342] + hash_xor_i[343] + hash_xor_i[344] + hash_xor_i[345] + hash_xor_i[346] + hash_xor_i[347] + hash_xor_i[348] + hash_xor_i[349] + hash_xor_i[350] + hash_xor_i[351] + hash_xor_i[352] + hash_xor_i[353] + hash_xor_i[354] + hash_xor_i[355] + hash_xor_i[356] + hash_xor_i[357] + hash_xor_i[358] + hash_xor_i[359] + hash_xor_i[360] + hash_xor_i[361] + hash_xor_i[362] + hash_xor_i[363] + hash_xor_i[364] + hash_xor_i[365] + hash_xor_i[366] + hash_xor_i[367] + hash_xor_i[368] + hash_xor_i[369] + hash_xor_i[370] + hash_xor_i[371] + hash_xor_i[372] + hash_xor_i[373] + hash_xor_i[374] + hash_xor_i[375] + hash_xor_i[376] + hash_xor_i[377] + hash_xor_i[378] + hash_xor_i[379] + hash_xor_i[380] + hash_xor_i[381] + hash_xor_i[382] + hash_xor_i[383] + hash_xor_i[384] + hash_xor_i[385] + hash_xor_i[386] + hash_xor_i[387] + hash_xor_i[388] + hash_xor_i[389] + hash_xor_i[390] + hash_xor_i[391] + hash_xor_i[392] + hash_xor_i[393] + hash_xor_i[394] + hash_xor_i[395] + hash_xor_i[396] + hash_xor_i[397] + hash_xor_i[398] + hash_xor_i[399] + hash_xor_i[400] + hash_xor_i[401] + hash_xor_i[402] + hash_xor_i[403] + hash_xor_i[404] + hash_xor_i[405] + hash_xor_i[406] + hash_xor_i[407] + hash_xor_i[408] + hash_xor_i[409] + hash_xor_i[410] + hash_xor_i[411] + hash_xor_i[412] + hash_xor_i[413] + hash_xor_i[414] + hash_xor_i[415] + hash_xor_i[416] + hash_xor_i[417] + hash_xor_i[418] + hash_xor_i[419] + hash_xor_i[420] + hash_xor_i[421] + hash_xor_i[422] + hash_xor_i[423] + hash_xor_i[424] + hash_xor_i[425] + hash_xor_i[426] + hash_xor_i[427] + hash_xor_i[428] + hash_xor_i[429] + hash_xor_i[430] + hash_xor_i[431] + hash_xor_i[432] + hash_xor_i[433] + hash_xor_i[434] + hash_xor_i[435] + hash_xor_i[436] + hash_xor_i[437] + hash_xor_i[438] + hash_xor_i[439] + hash_xor_i[440] + hash_xor_i[441] + hash_xor_i[442] + hash_xor_i[443] + hash_xor_i[444] + hash_xor_i[445] + hash_xor_i[446] + hash_xor_i[447] + hash_xor_i[448] + hash_xor_i[449] + hash_xor_i[450] + hash_xor_i[451] + hash_xor_i[452] + hash_xor_i[453] + hash_xor_i[454] + hash_xor_i[455] + hash_xor_i[456] + hash_xor_i[457] + hash_xor_i[458] + hash_xor_i[459] + hash_xor_i[460] + hash_xor_i[461] + hash_xor_i[462] + hash_xor_i[463] + hash_xor_i[464] + hash_xor_i[465] + hash_xor_i[466] + hash_xor_i[467] + hash_xor_i[468] + hash_xor_i[469] + hash_xor_i[470] + hash_xor_i[471] + hash_xor_i[472] + hash_xor_i[473] + hash_xor_i[474] + hash_xor_i[475] + hash_xor_i[476] + hash_xor_i[477] + hash_xor_i[478] + hash_xor_i[479] + hash_xor_i[480] + hash_xor_i[481] + hash_xor_i[482] + hash_xor_i[483] + hash_xor_i[484] + hash_xor_i[485] + hash_xor_i[486] + hash_xor_i[487] + hash_xor_i[488] + hash_xor_i[489] + hash_xor_i[490] + hash_xor_i[491] + hash_xor_i[492] + hash_xor_i[493] + hash_xor_i[494] + hash_xor_i[495] + hash_xor_i[496] + hash_xor_i[497] + hash_xor_i[498] + hash_xor_i[499] + hash_xor_i[500] + hash_xor_i[501] + hash_xor_i[502] + hash_xor_i[503] + hash_xor_i[504] + hash_xor_i[505] + hash_xor_i[506] + hash_xor_i[507] + hash_xor_i[508] + hash_xor_i[509] + hash_xor_i[510] + hash_xor_i[511] + hash_xor_i[512] + hash_xor_i[513] + hash_xor_i[514] + hash_xor_i[515] + hash_xor_i[516] + hash_xor_i[517] + hash_xor_i[518] + hash_xor_i[519] + hash_xor_i[520] + hash_xor_i[521] + hash_xor_i[522] + hash_xor_i[523] + hash_xor_i[524] + hash_xor_i[525] + hash_xor_i[526] + hash_xor_i[527] + hash_xor_i[528] + hash_xor_i[529] + hash_xor_i[530] + hash_xor_i[531] + hash_xor_i[532] + hash_xor_i[533] + hash_xor_i[534] + hash_xor_i[535] + hash_xor_i[536] + hash_xor_i[537] + hash_xor_i[538] + hash_xor_i[539] + hash_xor_i[540] + hash_xor_i[541] + hash_xor_i[542] + hash_xor_i[543] + hash_xor_i[544] + hash_xor_i[545] + hash_xor_i[546] + hash_xor_i[547] + hash_xor_i[548] + hash_xor_i[549] + hash_xor_i[550] + hash_xor_i[551] + hash_xor_i[552] + hash_xor_i[553] + hash_xor_i[554] + hash_xor_i[555] + hash_xor_i[556] + hash_xor_i[557] + hash_xor_i[558] + hash_xor_i[559] + hash_xor_i[560] + hash_xor_i[561] + hash_xor_i[562] + hash_xor_i[563] + hash_xor_i[564] + hash_xor_i[565] + hash_xor_i[566] + hash_xor_i[567] + hash_xor_i[568] + hash_xor_i[569] + hash_xor_i[570] + hash_xor_i[571] + hash_xor_i[572] + hash_xor_i[573] + hash_xor_i[574] + hash_xor_i[575] + hash_xor_i[576] + hash_xor_i[577] + hash_xor_i[578] + hash_xor_i[579] + hash_xor_i[580] + hash_xor_i[581] + hash_xor_i[582] + hash_xor_i[583] + hash_xor_i[584] + hash_xor_i[585] + hash_xor_i[586] + hash_xor_i[587] + hash_xor_i[588] + hash_xor_i[589] + hash_xor_i[590] + hash_xor_i[591] + hash_xor_i[592] + hash_xor_i[593] + hash_xor_i[594] + hash_xor_i[595] + hash_xor_i[596] + hash_xor_i[597] + hash_xor_i[598] + hash_xor_i[599] + hash_xor_i[600] + hash_xor_i[601] + hash_xor_i[602] + hash_xor_i[603] + hash_xor_i[604] + hash_xor_i[605] + hash_xor_i[606] + hash_xor_i[607] + hash_xor_i[608] + hash_xor_i[609] + hash_xor_i[610] + hash_xor_i[611] + hash_xor_i[612] + hash_xor_i[613] + hash_xor_i[614] + hash_xor_i[615] + hash_xor_i[616] + hash_xor_i[617] + hash_xor_i[618] + hash_xor_i[619] + hash_xor_i[620] + hash_xor_i[621] + hash_xor_i[622] + hash_xor_i[623] + hash_xor_i[624] + hash_xor_i[625] + hash_xor_i[626] + hash_xor_i[627] + hash_xor_i[628] + hash_xor_i[629] + hash_xor_i[630] + hash_xor_i[631] + hash_xor_i[632] + hash_xor_i[633] + hash_xor_i[634] + hash_xor_i[635] + hash_xor_i[636] + hash_xor_i[637] + hash_xor_i[638] + hash_xor_i[639] + hash_xor_i[640] + hash_xor_i[641] + hash_xor_i[642] + hash_xor_i[643] + hash_xor_i[644] + hash_xor_i[645] + hash_xor_i[646] + hash_xor_i[647] + hash_xor_i[648] + hash_xor_i[649] + hash_xor_i[650] + hash_xor_i[651] + hash_xor_i[652] + hash_xor_i[653] + hash_xor_i[654] + hash_xor_i[655] + hash_xor_i[656] + hash_xor_i[657] + hash_xor_i[658] + hash_xor_i[659] + hash_xor_i[660] + hash_xor_i[661] + hash_xor_i[662] + hash_xor_i[663] + hash_xor_i[664] + hash_xor_i[665] + hash_xor_i[666] + hash_xor_i[667] + hash_xor_i[668] + hash_xor_i[669] + hash_xor_i[670] + hash_xor_i[671] + hash_xor_i[672] + hash_xor_i[673] + hash_xor_i[674] + hash_xor_i[675] + hash_xor_i[676] + hash_xor_i[677] + hash_xor_i[678] + hash_xor_i[679] + hash_xor_i[680] + hash_xor_i[681] + hash_xor_i[682] + hash_xor_i[683] + hash_xor_i[684] + hash_xor_i[685] + hash_xor_i[686] + hash_xor_i[687] + hash_xor_i[688] + hash_xor_i[689] + hash_xor_i[690] + hash_xor_i[691] + hash_xor_i[692] + hash_xor_i[693] + hash_xor_i[694] + hash_xor_i[695] + hash_xor_i[696] + hash_xor_i[697] + hash_xor_i[698] + hash_xor_i[699] + hash_xor_i[700] + hash_xor_i[701] + hash_xor_i[702] + hash_xor_i[703] + hash_xor_i[704] + hash_xor_i[705] + hash_xor_i[706] + hash_xor_i[707] + hash_xor_i[708] + hash_xor_i[709] + hash_xor_i[710] + hash_xor_i[711] + hash_xor_i[712] + hash_xor_i[713] + hash_xor_i[714] + hash_xor_i[715] + hash_xor_i[716] + hash_xor_i[717] + hash_xor_i[718] + hash_xor_i[719] + hash_xor_i[720] + hash_xor_i[721] + hash_xor_i[722] + hash_xor_i[723] + hash_xor_i[724] + hash_xor_i[725] + hash_xor_i[726] + hash_xor_i[727] + hash_xor_i[728] + hash_xor_i[729] + hash_xor_i[730] + hash_xor_i[731] + hash_xor_i[732] + hash_xor_i[733] + hash_xor_i[734] + hash_xor_i[735] + hash_xor_i[736] + hash_xor_i[737] + hash_xor_i[738] + hash_xor_i[739] + hash_xor_i[740] + hash_xor_i[741] + hash_xor_i[742] + hash_xor_i[743] + hash_xor_i[744] + hash_xor_i[745] + hash_xor_i[746] + hash_xor_i[747] + hash_xor_i[748] + hash_xor_i[749] + hash_xor_i[750] + hash_xor_i[751] + hash_xor_i[752] + hash_xor_i[753] + hash_xor_i[754] + hash_xor_i[755] + hash_xor_i[756] + hash_xor_i[757] + hash_xor_i[758] + hash_xor_i[759] + hash_xor_i[760] + hash_xor_i[761] + hash_xor_i[762] + hash_xor_i[763] + hash_xor_i[764] + hash_xor_i[765] + hash_xor_i[766] + hash_xor_i[767] + hash_xor_i[768] + hash_xor_i[769] + hash_xor_i[770] + hash_xor_i[771] + hash_xor_i[772] + hash_xor_i[773] + hash_xor_i[774] + hash_xor_i[775] + hash_xor_i[776] + hash_xor_i[777] + hash_xor_i[778] + hash_xor_i[779] + hash_xor_i[780] + hash_xor_i[781] + hash_xor_i[782] + hash_xor_i[783] + hash_xor_i[784] + hash_xor_i[785] + hash_xor_i[786] + hash_xor_i[787] + hash_xor_i[788] + hash_xor_i[789] + hash_xor_i[790] + hash_xor_i[791] + hash_xor_i[792] + hash_xor_i[793] + hash_xor_i[794] + hash_xor_i[795] + hash_xor_i[796] + hash_xor_i[797] + hash_xor_i[798] + hash_xor_i[799] + hash_xor_i[800] + hash_xor_i[801] + hash_xor_i[802] + hash_xor_i[803] + hash_xor_i[804] + hash_xor_i[805] + hash_xor_i[806] + hash_xor_i[807] + hash_xor_i[808] + hash_xor_i[809] + hash_xor_i[810] + hash_xor_i[811] + hash_xor_i[812] + hash_xor_i[813] + hash_xor_i[814] + hash_xor_i[815] + hash_xor_i[816] + hash_xor_i[817] + hash_xor_i[818] + hash_xor_i[819] + hash_xor_i[820] + hash_xor_i[821] + hash_xor_i[822] + hash_xor_i[823] + hash_xor_i[824] + hash_xor_i[825] + hash_xor_i[826] + hash_xor_i[827] + hash_xor_i[828] + hash_xor_i[829] + hash_xor_i[830] + hash_xor_i[831] + hash_xor_i[832] + hash_xor_i[833] + hash_xor_i[834] + hash_xor_i[835] + hash_xor_i[836] + hash_xor_i[837] + hash_xor_i[838] + hash_xor_i[839] + hash_xor_i[840] + hash_xor_i[841] + hash_xor_i[842] + hash_xor_i[843] + hash_xor_i[844] + hash_xor_i[845] + hash_xor_i[846] + hash_xor_i[847] + hash_xor_i[848] + hash_xor_i[849] + hash_xor_i[850] + hash_xor_i[851] + hash_xor_i[852] + hash_xor_i[853] + hash_xor_i[854] + hash_xor_i[855] + hash_xor_i[856] + hash_xor_i[857] + hash_xor_i[858] + hash_xor_i[859] + hash_xor_i[860] + hash_xor_i[861] + hash_xor_i[862] + hash_xor_i[863] + hash_xor_i[864] + hash_xor_i[865] + hash_xor_i[866] + hash_xor_i[867] + hash_xor_i[868] + hash_xor_i[869] + hash_xor_i[870] + hash_xor_i[871] + hash_xor_i[872] + hash_xor_i[873] + hash_xor_i[874] + hash_xor_i[875] + hash_xor_i[876] + hash_xor_i[877] + hash_xor_i[878] + hash_xor_i[879] + hash_xor_i[880] + hash_xor_i[881] + hash_xor_i[882] + hash_xor_i[883] + hash_xor_i[884] + hash_xor_i[885] + hash_xor_i[886] + hash_xor_i[887] + hash_xor_i[888] + hash_xor_i[889] + hash_xor_i[890] + hash_xor_i[891] + hash_xor_i[892] + hash_xor_i[893] + hash_xor_i[894] + hash_xor_i[895] + hash_xor_i[896] + hash_xor_i[897] + hash_xor_i[898] + hash_xor_i[899] + hash_xor_i[900] + hash_xor_i[901] + hash_xor_i[902] + hash_xor_i[903] + hash_xor_i[904] + hash_xor_i[905] + hash_xor_i[906] + hash_xor_i[907] + hash_xor_i[908] + hash_xor_i[909] + hash_xor_i[910] + hash_xor_i[911] + hash_xor_i[912] + hash_xor_i[913] + hash_xor_i[914] + hash_xor_i[915] + hash_xor_i[916] + hash_xor_i[917] + hash_xor_i[918] + hash_xor_i[919] + hash_xor_i[920] + hash_xor_i[921] + hash_xor_i[922] + hash_xor_i[923] + hash_xor_i[924] + hash_xor_i[925] + hash_xor_i[926] + hash_xor_i[927] + hash_xor_i[928] + hash_xor_i[929] + hash_xor_i[930] + hash_xor_i[931] + hash_xor_i[932] + hash_xor_i[933] + hash_xor_i[934] + hash_xor_i[935] + hash_xor_i[936] + hash_xor_i[937] + hash_xor_i[938] + hash_xor_i[939] + hash_xor_i[940] + hash_xor_i[941] + hash_xor_i[942] + hash_xor_i[943] + hash_xor_i[944] + hash_xor_i[945] + hash_xor_i[946] + hash_xor_i[947] + hash_xor_i[948] + hash_xor_i[949] + hash_xor_i[950] + hash_xor_i[951] + hash_xor_i[952] + hash_xor_i[953] + hash_xor_i[954] + hash_xor_i[955] + hash_xor_i[956] + hash_xor_i[957] + hash_xor_i[958] + hash_xor_i[959] + hash_xor_i[960] + hash_xor_i[961] + hash_xor_i[962] + hash_xor_i[963] + hash_xor_i[964] + hash_xor_i[965] + hash_xor_i[966] + hash_xor_i[967] + hash_xor_i[968] + hash_xor_i[969] + hash_xor_i[970] + hash_xor_i[971] + hash_xor_i[972] + hash_xor_i[973] + hash_xor_i[974] + hash_xor_i[975] + hash_xor_i[976] + hash_xor_i[977] + hash_xor_i[978] + hash_xor_i[979] + hash_xor_i[980] + hash_xor_i[981] + hash_xor_i[982] + hash_xor_i[983] + hash_xor_i[984] + hash_xor_i[985] + hash_xor_i[986] + hash_xor_i[987] + hash_xor_i[988] + hash_xor_i[989] + hash_xor_i[990] + hash_xor_i[991] + hash_xor_i[992] + hash_xor_i[993] + hash_xor_i[994] + hash_xor_i[995] + hash_xor_i[996] + hash_xor_i[997] + hash_xor_i[998] + hash_xor_i[999] + hash_xor_i[1000] + hash_xor_i[1001] + hash_xor_i[1002] + hash_xor_i[1003] + hash_xor_i[1004] + hash_xor_i[1005] + hash_xor_i[1006] + hash_xor_i[1007] + hash_xor_i[1008] + hash_xor_i[1009] + hash_xor_i[1010] + hash_xor_i[1011] + hash_xor_i[1012] + hash_xor_i[1013] + hash_xor_i[1014] + hash_xor_i[1015] + hash_xor_i[1016] + hash_xor_i[1017] + hash_xor_i[1018] + hash_xor_i[1019] + hash_xor_i[1020] + hash_xor_i[1021] + hash_xor_i[1022] + hash_xor_i[1023];

end

endmodule
