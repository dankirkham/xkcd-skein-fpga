module input_register (
	input clk_i,
	input rst_i,
	input [1023:0] output_register_i,
	output 
	
endmodule