module header_constant (
  output [7:0] output_o
);

assign output_o = 8'h9A;

endmodule
