// TODO: This module is not currently used. It will probably synthesize faster.
// To use this it, it must be verified with block_ram_test. It has already been
// verified with Verilator.

module block_ram_multidimensional (
  input clk_i,
  input write_i,
  input [15:0] data_i,
  input [7:0] address_i,

  output reg [15:0] data_o
);

reg [15:0] data_d [255:0];
reg [15:0] data_q [255:0];

// Read Mux
always @(*) begin
  data_o = data_q[address_i];
end

// Write mux - generated by ./gen/write_mux_multidimensional.py
always @(*) begin
  if (write_i == 1'b1) begin
    if (address_i == 8'd0) begin
      data_d[0] = data_i;
      data_d[255:1] = data_q[255:1];
    end else if (address_i == 8'd1) begin
      data_d[0] = data_q[0];
      data_d[1] = data_i;
      data_d[255:2] = data_q[255:2];
    end else if (address_i == 8'd2) begin
      data_d[1:0] = data_q[1:0];
      data_d[2] = data_i;
      data_d[255:3] = data_q[255:3];
    end else if (address_i == 8'd3) begin
      data_d[2:0] = data_q[2:0];
      data_d[3] = data_i;
      data_d[255:4] = data_q[255:4];
    end else if (address_i == 8'd4) begin
      data_d[3:0] = data_q[3:0];
      data_d[4] = data_i;
      data_d[255:5] = data_q[255:5];
    end else if (address_i == 8'd5) begin
      data_d[4:0] = data_q[4:0];
      data_d[5] = data_i;
      data_d[255:6] = data_q[255:6];
    end else if (address_i == 8'd6) begin
      data_d[5:0] = data_q[5:0];
      data_d[6] = data_i;
      data_d[255:7] = data_q[255:7];
    end else if (address_i == 8'd7) begin
      data_d[6:0] = data_q[6:0];
      data_d[7] = data_i;
      data_d[255:8] = data_q[255:8];
    end else if (address_i == 8'd8) begin
      data_d[7:0] = data_q[7:0];
      data_d[8] = data_i;
      data_d[255:9] = data_q[255:9];
    end else if (address_i == 8'd9) begin
      data_d[8:0] = data_q[8:0];
      data_d[9] = data_i;
      data_d[255:10] = data_q[255:10];
    end else if (address_i == 8'd10) begin
      data_d[9:0] = data_q[9:0];
      data_d[10] = data_i;
      data_d[255:11] = data_q[255:11];
    end else if (address_i == 8'd11) begin
      data_d[10:0] = data_q[10:0];
      data_d[11] = data_i;
      data_d[255:12] = data_q[255:12];
    end else if (address_i == 8'd12) begin
      data_d[11:0] = data_q[11:0];
      data_d[12] = data_i;
      data_d[255:13] = data_q[255:13];
    end else if (address_i == 8'd13) begin
      data_d[12:0] = data_q[12:0];
      data_d[13] = data_i;
      data_d[255:14] = data_q[255:14];
    end else if (address_i == 8'd14) begin
      data_d[13:0] = data_q[13:0];
      data_d[14] = data_i;
      data_d[255:15] = data_q[255:15];
    end else if (address_i == 8'd15) begin
      data_d[14:0] = data_q[14:0];
      data_d[15] = data_i;
      data_d[255:16] = data_q[255:16];
    end else if (address_i == 8'd16) begin
      data_d[15:0] = data_q[15:0];
      data_d[16] = data_i;
      data_d[255:17] = data_q[255:17];
    end else if (address_i == 8'd17) begin
      data_d[16:0] = data_q[16:0];
      data_d[17] = data_i;
      data_d[255:18] = data_q[255:18];
    end else if (address_i == 8'd18) begin
      data_d[17:0] = data_q[17:0];
      data_d[18] = data_i;
      data_d[255:19] = data_q[255:19];
    end else if (address_i == 8'd19) begin
      data_d[18:0] = data_q[18:0];
      data_d[19] = data_i;
      data_d[255:20] = data_q[255:20];
    end else if (address_i == 8'd20) begin
      data_d[19:0] = data_q[19:0];
      data_d[20] = data_i;
      data_d[255:21] = data_q[255:21];
    end else if (address_i == 8'd21) begin
      data_d[20:0] = data_q[20:0];
      data_d[21] = data_i;
      data_d[255:22] = data_q[255:22];
    end else if (address_i == 8'd22) begin
      data_d[21:0] = data_q[21:0];
      data_d[22] = data_i;
      data_d[255:23] = data_q[255:23];
    end else if (address_i == 8'd23) begin
      data_d[22:0] = data_q[22:0];
      data_d[23] = data_i;
      data_d[255:24] = data_q[255:24];
    end else if (address_i == 8'd24) begin
      data_d[23:0] = data_q[23:0];
      data_d[24] = data_i;
      data_d[255:25] = data_q[255:25];
    end else if (address_i == 8'd25) begin
      data_d[24:0] = data_q[24:0];
      data_d[25] = data_i;
      data_d[255:26] = data_q[255:26];
    end else if (address_i == 8'd26) begin
      data_d[25:0] = data_q[25:0];
      data_d[26] = data_i;
      data_d[255:27] = data_q[255:27];
    end else if (address_i == 8'd27) begin
      data_d[26:0] = data_q[26:0];
      data_d[27] = data_i;
      data_d[255:28] = data_q[255:28];
    end else if (address_i == 8'd28) begin
      data_d[27:0] = data_q[27:0];
      data_d[28] = data_i;
      data_d[255:29] = data_q[255:29];
    end else if (address_i == 8'd29) begin
      data_d[28:0] = data_q[28:0];
      data_d[29] = data_i;
      data_d[255:30] = data_q[255:30];
    end else if (address_i == 8'd30) begin
      data_d[29:0] = data_q[29:0];
      data_d[30] = data_i;
      data_d[255:31] = data_q[255:31];
    end else if (address_i == 8'd31) begin
      data_d[30:0] = data_q[30:0];
      data_d[31] = data_i;
      data_d[255:32] = data_q[255:32];
    end else if (address_i == 8'd32) begin
      data_d[31:0] = data_q[31:0];
      data_d[32] = data_i;
      data_d[255:33] = data_q[255:33];
    end else if (address_i == 8'd33) begin
      data_d[32:0] = data_q[32:0];
      data_d[33] = data_i;
      data_d[255:34] = data_q[255:34];
    end else if (address_i == 8'd34) begin
      data_d[33:0] = data_q[33:0];
      data_d[34] = data_i;
      data_d[255:35] = data_q[255:35];
    end else if (address_i == 8'd35) begin
      data_d[34:0] = data_q[34:0];
      data_d[35] = data_i;
      data_d[255:36] = data_q[255:36];
    end else if (address_i == 8'd36) begin
      data_d[35:0] = data_q[35:0];
      data_d[36] = data_i;
      data_d[255:37] = data_q[255:37];
    end else if (address_i == 8'd37) begin
      data_d[36:0] = data_q[36:0];
      data_d[37] = data_i;
      data_d[255:38] = data_q[255:38];
    end else if (address_i == 8'd38) begin
      data_d[37:0] = data_q[37:0];
      data_d[38] = data_i;
      data_d[255:39] = data_q[255:39];
    end else if (address_i == 8'd39) begin
      data_d[38:0] = data_q[38:0];
      data_d[39] = data_i;
      data_d[255:40] = data_q[255:40];
    end else if (address_i == 8'd40) begin
      data_d[39:0] = data_q[39:0];
      data_d[40] = data_i;
      data_d[255:41] = data_q[255:41];
    end else if (address_i == 8'd41) begin
      data_d[40:0] = data_q[40:0];
      data_d[41] = data_i;
      data_d[255:42] = data_q[255:42];
    end else if (address_i == 8'd42) begin
      data_d[41:0] = data_q[41:0];
      data_d[42] = data_i;
      data_d[255:43] = data_q[255:43];
    end else if (address_i == 8'd43) begin
      data_d[42:0] = data_q[42:0];
      data_d[43] = data_i;
      data_d[255:44] = data_q[255:44];
    end else if (address_i == 8'd44) begin
      data_d[43:0] = data_q[43:0];
      data_d[44] = data_i;
      data_d[255:45] = data_q[255:45];
    end else if (address_i == 8'd45) begin
      data_d[44:0] = data_q[44:0];
      data_d[45] = data_i;
      data_d[255:46] = data_q[255:46];
    end else if (address_i == 8'd46) begin
      data_d[45:0] = data_q[45:0];
      data_d[46] = data_i;
      data_d[255:47] = data_q[255:47];
    end else if (address_i == 8'd47) begin
      data_d[46:0] = data_q[46:0];
      data_d[47] = data_i;
      data_d[255:48] = data_q[255:48];
    end else if (address_i == 8'd48) begin
      data_d[47:0] = data_q[47:0];
      data_d[48] = data_i;
      data_d[255:49] = data_q[255:49];
    end else if (address_i == 8'd49) begin
      data_d[48:0] = data_q[48:0];
      data_d[49] = data_i;
      data_d[255:50] = data_q[255:50];
    end else if (address_i == 8'd50) begin
      data_d[49:0] = data_q[49:0];
      data_d[50] = data_i;
      data_d[255:51] = data_q[255:51];
    end else if (address_i == 8'd51) begin
      data_d[50:0] = data_q[50:0];
      data_d[51] = data_i;
      data_d[255:52] = data_q[255:52];
    end else if (address_i == 8'd52) begin
      data_d[51:0] = data_q[51:0];
      data_d[52] = data_i;
      data_d[255:53] = data_q[255:53];
    end else if (address_i == 8'd53) begin
      data_d[52:0] = data_q[52:0];
      data_d[53] = data_i;
      data_d[255:54] = data_q[255:54];
    end else if (address_i == 8'd54) begin
      data_d[53:0] = data_q[53:0];
      data_d[54] = data_i;
      data_d[255:55] = data_q[255:55];
    end else if (address_i == 8'd55) begin
      data_d[54:0] = data_q[54:0];
      data_d[55] = data_i;
      data_d[255:56] = data_q[255:56];
    end else if (address_i == 8'd56) begin
      data_d[55:0] = data_q[55:0];
      data_d[56] = data_i;
      data_d[255:57] = data_q[255:57];
    end else if (address_i == 8'd57) begin
      data_d[56:0] = data_q[56:0];
      data_d[57] = data_i;
      data_d[255:58] = data_q[255:58];
    end else if (address_i == 8'd58) begin
      data_d[57:0] = data_q[57:0];
      data_d[58] = data_i;
      data_d[255:59] = data_q[255:59];
    end else if (address_i == 8'd59) begin
      data_d[58:0] = data_q[58:0];
      data_d[59] = data_i;
      data_d[255:60] = data_q[255:60];
    end else if (address_i == 8'd60) begin
      data_d[59:0] = data_q[59:0];
      data_d[60] = data_i;
      data_d[255:61] = data_q[255:61];
    end else if (address_i == 8'd61) begin
      data_d[60:0] = data_q[60:0];
      data_d[61] = data_i;
      data_d[255:62] = data_q[255:62];
    end else if (address_i == 8'd62) begin
      data_d[61:0] = data_q[61:0];
      data_d[62] = data_i;
      data_d[255:63] = data_q[255:63];
    end else if (address_i == 8'd63) begin
      data_d[62:0] = data_q[62:0];
      data_d[63] = data_i;
      data_d[255:64] = data_q[255:64];
    end else if (address_i == 8'd64) begin
      data_d[63:0] = data_q[63:0];
      data_d[64] = data_i;
      data_d[255:65] = data_q[255:65];
    end else if (address_i == 8'd65) begin
      data_d[64:0] = data_q[64:0];
      data_d[65] = data_i;
      data_d[255:66] = data_q[255:66];
    end else if (address_i == 8'd66) begin
      data_d[65:0] = data_q[65:0];
      data_d[66] = data_i;
      data_d[255:67] = data_q[255:67];
    end else if (address_i == 8'd67) begin
      data_d[66:0] = data_q[66:0];
      data_d[67] = data_i;
      data_d[255:68] = data_q[255:68];
    end else if (address_i == 8'd68) begin
      data_d[67:0] = data_q[67:0];
      data_d[68] = data_i;
      data_d[255:69] = data_q[255:69];
    end else if (address_i == 8'd69) begin
      data_d[68:0] = data_q[68:0];
      data_d[69] = data_i;
      data_d[255:70] = data_q[255:70];
    end else if (address_i == 8'd70) begin
      data_d[69:0] = data_q[69:0];
      data_d[70] = data_i;
      data_d[255:71] = data_q[255:71];
    end else if (address_i == 8'd71) begin
      data_d[70:0] = data_q[70:0];
      data_d[71] = data_i;
      data_d[255:72] = data_q[255:72];
    end else if (address_i == 8'd72) begin
      data_d[71:0] = data_q[71:0];
      data_d[72] = data_i;
      data_d[255:73] = data_q[255:73];
    end else if (address_i == 8'd73) begin
      data_d[72:0] = data_q[72:0];
      data_d[73] = data_i;
      data_d[255:74] = data_q[255:74];
    end else if (address_i == 8'd74) begin
      data_d[73:0] = data_q[73:0];
      data_d[74] = data_i;
      data_d[255:75] = data_q[255:75];
    end else if (address_i == 8'd75) begin
      data_d[74:0] = data_q[74:0];
      data_d[75] = data_i;
      data_d[255:76] = data_q[255:76];
    end else if (address_i == 8'd76) begin
      data_d[75:0] = data_q[75:0];
      data_d[76] = data_i;
      data_d[255:77] = data_q[255:77];
    end else if (address_i == 8'd77) begin
      data_d[76:0] = data_q[76:0];
      data_d[77] = data_i;
      data_d[255:78] = data_q[255:78];
    end else if (address_i == 8'd78) begin
      data_d[77:0] = data_q[77:0];
      data_d[78] = data_i;
      data_d[255:79] = data_q[255:79];
    end else if (address_i == 8'd79) begin
      data_d[78:0] = data_q[78:0];
      data_d[79] = data_i;
      data_d[255:80] = data_q[255:80];
    end else if (address_i == 8'd80) begin
      data_d[79:0] = data_q[79:0];
      data_d[80] = data_i;
      data_d[255:81] = data_q[255:81];
    end else if (address_i == 8'd81) begin
      data_d[80:0] = data_q[80:0];
      data_d[81] = data_i;
      data_d[255:82] = data_q[255:82];
    end else if (address_i == 8'd82) begin
      data_d[81:0] = data_q[81:0];
      data_d[82] = data_i;
      data_d[255:83] = data_q[255:83];
    end else if (address_i == 8'd83) begin
      data_d[82:0] = data_q[82:0];
      data_d[83] = data_i;
      data_d[255:84] = data_q[255:84];
    end else if (address_i == 8'd84) begin
      data_d[83:0] = data_q[83:0];
      data_d[84] = data_i;
      data_d[255:85] = data_q[255:85];
    end else if (address_i == 8'd85) begin
      data_d[84:0] = data_q[84:0];
      data_d[85] = data_i;
      data_d[255:86] = data_q[255:86];
    end else if (address_i == 8'd86) begin
      data_d[85:0] = data_q[85:0];
      data_d[86] = data_i;
      data_d[255:87] = data_q[255:87];
    end else if (address_i == 8'd87) begin
      data_d[86:0] = data_q[86:0];
      data_d[87] = data_i;
      data_d[255:88] = data_q[255:88];
    end else if (address_i == 8'd88) begin
      data_d[87:0] = data_q[87:0];
      data_d[88] = data_i;
      data_d[255:89] = data_q[255:89];
    end else if (address_i == 8'd89) begin
      data_d[88:0] = data_q[88:0];
      data_d[89] = data_i;
      data_d[255:90] = data_q[255:90];
    end else if (address_i == 8'd90) begin
      data_d[89:0] = data_q[89:0];
      data_d[90] = data_i;
      data_d[255:91] = data_q[255:91];
    end else if (address_i == 8'd91) begin
      data_d[90:0] = data_q[90:0];
      data_d[91] = data_i;
      data_d[255:92] = data_q[255:92];
    end else if (address_i == 8'd92) begin
      data_d[91:0] = data_q[91:0];
      data_d[92] = data_i;
      data_d[255:93] = data_q[255:93];
    end else if (address_i == 8'd93) begin
      data_d[92:0] = data_q[92:0];
      data_d[93] = data_i;
      data_d[255:94] = data_q[255:94];
    end else if (address_i == 8'd94) begin
      data_d[93:0] = data_q[93:0];
      data_d[94] = data_i;
      data_d[255:95] = data_q[255:95];
    end else if (address_i == 8'd95) begin
      data_d[94:0] = data_q[94:0];
      data_d[95] = data_i;
      data_d[255:96] = data_q[255:96];
    end else if (address_i == 8'd96) begin
      data_d[95:0] = data_q[95:0];
      data_d[96] = data_i;
      data_d[255:97] = data_q[255:97];
    end else if (address_i == 8'd97) begin
      data_d[96:0] = data_q[96:0];
      data_d[97] = data_i;
      data_d[255:98] = data_q[255:98];
    end else if (address_i == 8'd98) begin
      data_d[97:0] = data_q[97:0];
      data_d[98] = data_i;
      data_d[255:99] = data_q[255:99];
    end else if (address_i == 8'd99) begin
      data_d[98:0] = data_q[98:0];
      data_d[99] = data_i;
      data_d[255:100] = data_q[255:100];
    end else if (address_i == 8'd100) begin
      data_d[99:0] = data_q[99:0];
      data_d[100] = data_i;
      data_d[255:101] = data_q[255:101];
    end else if (address_i == 8'd101) begin
      data_d[100:0] = data_q[100:0];
      data_d[101] = data_i;
      data_d[255:102] = data_q[255:102];
    end else if (address_i == 8'd102) begin
      data_d[101:0] = data_q[101:0];
      data_d[102] = data_i;
      data_d[255:103] = data_q[255:103];
    end else if (address_i == 8'd103) begin
      data_d[102:0] = data_q[102:0];
      data_d[103] = data_i;
      data_d[255:104] = data_q[255:104];
    end else if (address_i == 8'd104) begin
      data_d[103:0] = data_q[103:0];
      data_d[104] = data_i;
      data_d[255:105] = data_q[255:105];
    end else if (address_i == 8'd105) begin
      data_d[104:0] = data_q[104:0];
      data_d[105] = data_i;
      data_d[255:106] = data_q[255:106];
    end else if (address_i == 8'd106) begin
      data_d[105:0] = data_q[105:0];
      data_d[106] = data_i;
      data_d[255:107] = data_q[255:107];
    end else if (address_i == 8'd107) begin
      data_d[106:0] = data_q[106:0];
      data_d[107] = data_i;
      data_d[255:108] = data_q[255:108];
    end else if (address_i == 8'd108) begin
      data_d[107:0] = data_q[107:0];
      data_d[108] = data_i;
      data_d[255:109] = data_q[255:109];
    end else if (address_i == 8'd109) begin
      data_d[108:0] = data_q[108:0];
      data_d[109] = data_i;
      data_d[255:110] = data_q[255:110];
    end else if (address_i == 8'd110) begin
      data_d[109:0] = data_q[109:0];
      data_d[110] = data_i;
      data_d[255:111] = data_q[255:111];
    end else if (address_i == 8'd111) begin
      data_d[110:0] = data_q[110:0];
      data_d[111] = data_i;
      data_d[255:112] = data_q[255:112];
    end else if (address_i == 8'd112) begin
      data_d[111:0] = data_q[111:0];
      data_d[112] = data_i;
      data_d[255:113] = data_q[255:113];
    end else if (address_i == 8'd113) begin
      data_d[112:0] = data_q[112:0];
      data_d[113] = data_i;
      data_d[255:114] = data_q[255:114];
    end else if (address_i == 8'd114) begin
      data_d[113:0] = data_q[113:0];
      data_d[114] = data_i;
      data_d[255:115] = data_q[255:115];
    end else if (address_i == 8'd115) begin
      data_d[114:0] = data_q[114:0];
      data_d[115] = data_i;
      data_d[255:116] = data_q[255:116];
    end else if (address_i == 8'd116) begin
      data_d[115:0] = data_q[115:0];
      data_d[116] = data_i;
      data_d[255:117] = data_q[255:117];
    end else if (address_i == 8'd117) begin
      data_d[116:0] = data_q[116:0];
      data_d[117] = data_i;
      data_d[255:118] = data_q[255:118];
    end else if (address_i == 8'd118) begin
      data_d[117:0] = data_q[117:0];
      data_d[118] = data_i;
      data_d[255:119] = data_q[255:119];
    end else if (address_i == 8'd119) begin
      data_d[118:0] = data_q[118:0];
      data_d[119] = data_i;
      data_d[255:120] = data_q[255:120];
    end else if (address_i == 8'd120) begin
      data_d[119:0] = data_q[119:0];
      data_d[120] = data_i;
      data_d[255:121] = data_q[255:121];
    end else if (address_i == 8'd121) begin
      data_d[120:0] = data_q[120:0];
      data_d[121] = data_i;
      data_d[255:122] = data_q[255:122];
    end else if (address_i == 8'd122) begin
      data_d[121:0] = data_q[121:0];
      data_d[122] = data_i;
      data_d[255:123] = data_q[255:123];
    end else if (address_i == 8'd123) begin
      data_d[122:0] = data_q[122:0];
      data_d[123] = data_i;
      data_d[255:124] = data_q[255:124];
    end else if (address_i == 8'd124) begin
      data_d[123:0] = data_q[123:0];
      data_d[124] = data_i;
      data_d[255:125] = data_q[255:125];
    end else if (address_i == 8'd125) begin
      data_d[124:0] = data_q[124:0];
      data_d[125] = data_i;
      data_d[255:126] = data_q[255:126];
    end else if (address_i == 8'd126) begin
      data_d[125:0] = data_q[125:0];
      data_d[126] = data_i;
      data_d[255:127] = data_q[255:127];
    end else if (address_i == 8'd127) begin
      data_d[126:0] = data_q[126:0];
      data_d[127] = data_i;
      data_d[255:128] = data_q[255:128];
    end else if (address_i == 8'd128) begin
      data_d[127:0] = data_q[127:0];
      data_d[128] = data_i;
      data_d[255:129] = data_q[255:129];
    end else if (address_i == 8'd129) begin
      data_d[128:0] = data_q[128:0];
      data_d[129] = data_i;
      data_d[255:130] = data_q[255:130];
    end else if (address_i == 8'd130) begin
      data_d[129:0] = data_q[129:0];
      data_d[130] = data_i;
      data_d[255:131] = data_q[255:131];
    end else if (address_i == 8'd131) begin
      data_d[130:0] = data_q[130:0];
      data_d[131] = data_i;
      data_d[255:132] = data_q[255:132];
    end else if (address_i == 8'd132) begin
      data_d[131:0] = data_q[131:0];
      data_d[132] = data_i;
      data_d[255:133] = data_q[255:133];
    end else if (address_i == 8'd133) begin
      data_d[132:0] = data_q[132:0];
      data_d[133] = data_i;
      data_d[255:134] = data_q[255:134];
    end else if (address_i == 8'd134) begin
      data_d[133:0] = data_q[133:0];
      data_d[134] = data_i;
      data_d[255:135] = data_q[255:135];
    end else if (address_i == 8'd135) begin
      data_d[134:0] = data_q[134:0];
      data_d[135] = data_i;
      data_d[255:136] = data_q[255:136];
    end else if (address_i == 8'd136) begin
      data_d[135:0] = data_q[135:0];
      data_d[136] = data_i;
      data_d[255:137] = data_q[255:137];
    end else if (address_i == 8'd137) begin
      data_d[136:0] = data_q[136:0];
      data_d[137] = data_i;
      data_d[255:138] = data_q[255:138];
    end else if (address_i == 8'd138) begin
      data_d[137:0] = data_q[137:0];
      data_d[138] = data_i;
      data_d[255:139] = data_q[255:139];
    end else if (address_i == 8'd139) begin
      data_d[138:0] = data_q[138:0];
      data_d[139] = data_i;
      data_d[255:140] = data_q[255:140];
    end else if (address_i == 8'd140) begin
      data_d[139:0] = data_q[139:0];
      data_d[140] = data_i;
      data_d[255:141] = data_q[255:141];
    end else if (address_i == 8'd141) begin
      data_d[140:0] = data_q[140:0];
      data_d[141] = data_i;
      data_d[255:142] = data_q[255:142];
    end else if (address_i == 8'd142) begin
      data_d[141:0] = data_q[141:0];
      data_d[142] = data_i;
      data_d[255:143] = data_q[255:143];
    end else if (address_i == 8'd143) begin
      data_d[142:0] = data_q[142:0];
      data_d[143] = data_i;
      data_d[255:144] = data_q[255:144];
    end else if (address_i == 8'd144) begin
      data_d[143:0] = data_q[143:0];
      data_d[144] = data_i;
      data_d[255:145] = data_q[255:145];
    end else if (address_i == 8'd145) begin
      data_d[144:0] = data_q[144:0];
      data_d[145] = data_i;
      data_d[255:146] = data_q[255:146];
    end else if (address_i == 8'd146) begin
      data_d[145:0] = data_q[145:0];
      data_d[146] = data_i;
      data_d[255:147] = data_q[255:147];
    end else if (address_i == 8'd147) begin
      data_d[146:0] = data_q[146:0];
      data_d[147] = data_i;
      data_d[255:148] = data_q[255:148];
    end else if (address_i == 8'd148) begin
      data_d[147:0] = data_q[147:0];
      data_d[148] = data_i;
      data_d[255:149] = data_q[255:149];
    end else if (address_i == 8'd149) begin
      data_d[148:0] = data_q[148:0];
      data_d[149] = data_i;
      data_d[255:150] = data_q[255:150];
    end else if (address_i == 8'd150) begin
      data_d[149:0] = data_q[149:0];
      data_d[150] = data_i;
      data_d[255:151] = data_q[255:151];
    end else if (address_i == 8'd151) begin
      data_d[150:0] = data_q[150:0];
      data_d[151] = data_i;
      data_d[255:152] = data_q[255:152];
    end else if (address_i == 8'd152) begin
      data_d[151:0] = data_q[151:0];
      data_d[152] = data_i;
      data_d[255:153] = data_q[255:153];
    end else if (address_i == 8'd153) begin
      data_d[152:0] = data_q[152:0];
      data_d[153] = data_i;
      data_d[255:154] = data_q[255:154];
    end else if (address_i == 8'd154) begin
      data_d[153:0] = data_q[153:0];
      data_d[154] = data_i;
      data_d[255:155] = data_q[255:155];
    end else if (address_i == 8'd155) begin
      data_d[154:0] = data_q[154:0];
      data_d[155] = data_i;
      data_d[255:156] = data_q[255:156];
    end else if (address_i == 8'd156) begin
      data_d[155:0] = data_q[155:0];
      data_d[156] = data_i;
      data_d[255:157] = data_q[255:157];
    end else if (address_i == 8'd157) begin
      data_d[156:0] = data_q[156:0];
      data_d[157] = data_i;
      data_d[255:158] = data_q[255:158];
    end else if (address_i == 8'd158) begin
      data_d[157:0] = data_q[157:0];
      data_d[158] = data_i;
      data_d[255:159] = data_q[255:159];
    end else if (address_i == 8'd159) begin
      data_d[158:0] = data_q[158:0];
      data_d[159] = data_i;
      data_d[255:160] = data_q[255:160];
    end else if (address_i == 8'd160) begin
      data_d[159:0] = data_q[159:0];
      data_d[160] = data_i;
      data_d[255:161] = data_q[255:161];
    end else if (address_i == 8'd161) begin
      data_d[160:0] = data_q[160:0];
      data_d[161] = data_i;
      data_d[255:162] = data_q[255:162];
    end else if (address_i == 8'd162) begin
      data_d[161:0] = data_q[161:0];
      data_d[162] = data_i;
      data_d[255:163] = data_q[255:163];
    end else if (address_i == 8'd163) begin
      data_d[162:0] = data_q[162:0];
      data_d[163] = data_i;
      data_d[255:164] = data_q[255:164];
    end else if (address_i == 8'd164) begin
      data_d[163:0] = data_q[163:0];
      data_d[164] = data_i;
      data_d[255:165] = data_q[255:165];
    end else if (address_i == 8'd165) begin
      data_d[164:0] = data_q[164:0];
      data_d[165] = data_i;
      data_d[255:166] = data_q[255:166];
    end else if (address_i == 8'd166) begin
      data_d[165:0] = data_q[165:0];
      data_d[166] = data_i;
      data_d[255:167] = data_q[255:167];
    end else if (address_i == 8'd167) begin
      data_d[166:0] = data_q[166:0];
      data_d[167] = data_i;
      data_d[255:168] = data_q[255:168];
    end else if (address_i == 8'd168) begin
      data_d[167:0] = data_q[167:0];
      data_d[168] = data_i;
      data_d[255:169] = data_q[255:169];
    end else if (address_i == 8'd169) begin
      data_d[168:0] = data_q[168:0];
      data_d[169] = data_i;
      data_d[255:170] = data_q[255:170];
    end else if (address_i == 8'd170) begin
      data_d[169:0] = data_q[169:0];
      data_d[170] = data_i;
      data_d[255:171] = data_q[255:171];
    end else if (address_i == 8'd171) begin
      data_d[170:0] = data_q[170:0];
      data_d[171] = data_i;
      data_d[255:172] = data_q[255:172];
    end else if (address_i == 8'd172) begin
      data_d[171:0] = data_q[171:0];
      data_d[172] = data_i;
      data_d[255:173] = data_q[255:173];
    end else if (address_i == 8'd173) begin
      data_d[172:0] = data_q[172:0];
      data_d[173] = data_i;
      data_d[255:174] = data_q[255:174];
    end else if (address_i == 8'd174) begin
      data_d[173:0] = data_q[173:0];
      data_d[174] = data_i;
      data_d[255:175] = data_q[255:175];
    end else if (address_i == 8'd175) begin
      data_d[174:0] = data_q[174:0];
      data_d[175] = data_i;
      data_d[255:176] = data_q[255:176];
    end else if (address_i == 8'd176) begin
      data_d[175:0] = data_q[175:0];
      data_d[176] = data_i;
      data_d[255:177] = data_q[255:177];
    end else if (address_i == 8'd177) begin
      data_d[176:0] = data_q[176:0];
      data_d[177] = data_i;
      data_d[255:178] = data_q[255:178];
    end else if (address_i == 8'd178) begin
      data_d[177:0] = data_q[177:0];
      data_d[178] = data_i;
      data_d[255:179] = data_q[255:179];
    end else if (address_i == 8'd179) begin
      data_d[178:0] = data_q[178:0];
      data_d[179] = data_i;
      data_d[255:180] = data_q[255:180];
    end else if (address_i == 8'd180) begin
      data_d[179:0] = data_q[179:0];
      data_d[180] = data_i;
      data_d[255:181] = data_q[255:181];
    end else if (address_i == 8'd181) begin
      data_d[180:0] = data_q[180:0];
      data_d[181] = data_i;
      data_d[255:182] = data_q[255:182];
    end else if (address_i == 8'd182) begin
      data_d[181:0] = data_q[181:0];
      data_d[182] = data_i;
      data_d[255:183] = data_q[255:183];
    end else if (address_i == 8'd183) begin
      data_d[182:0] = data_q[182:0];
      data_d[183] = data_i;
      data_d[255:184] = data_q[255:184];
    end else if (address_i == 8'd184) begin
      data_d[183:0] = data_q[183:0];
      data_d[184] = data_i;
      data_d[255:185] = data_q[255:185];
    end else if (address_i == 8'd185) begin
      data_d[184:0] = data_q[184:0];
      data_d[185] = data_i;
      data_d[255:186] = data_q[255:186];
    end else if (address_i == 8'd186) begin
      data_d[185:0] = data_q[185:0];
      data_d[186] = data_i;
      data_d[255:187] = data_q[255:187];
    end else if (address_i == 8'd187) begin
      data_d[186:0] = data_q[186:0];
      data_d[187] = data_i;
      data_d[255:188] = data_q[255:188];
    end else if (address_i == 8'd188) begin
      data_d[187:0] = data_q[187:0];
      data_d[188] = data_i;
      data_d[255:189] = data_q[255:189];
    end else if (address_i == 8'd189) begin
      data_d[188:0] = data_q[188:0];
      data_d[189] = data_i;
      data_d[255:190] = data_q[255:190];
    end else if (address_i == 8'd190) begin
      data_d[189:0] = data_q[189:0];
      data_d[190] = data_i;
      data_d[255:191] = data_q[255:191];
    end else if (address_i == 8'd191) begin
      data_d[190:0] = data_q[190:0];
      data_d[191] = data_i;
      data_d[255:192] = data_q[255:192];
    end else if (address_i == 8'd192) begin
      data_d[191:0] = data_q[191:0];
      data_d[192] = data_i;
      data_d[255:193] = data_q[255:193];
    end else if (address_i == 8'd193) begin
      data_d[192:0] = data_q[192:0];
      data_d[193] = data_i;
      data_d[255:194] = data_q[255:194];
    end else if (address_i == 8'd194) begin
      data_d[193:0] = data_q[193:0];
      data_d[194] = data_i;
      data_d[255:195] = data_q[255:195];
    end else if (address_i == 8'd195) begin
      data_d[194:0] = data_q[194:0];
      data_d[195] = data_i;
      data_d[255:196] = data_q[255:196];
    end else if (address_i == 8'd196) begin
      data_d[195:0] = data_q[195:0];
      data_d[196] = data_i;
      data_d[255:197] = data_q[255:197];
    end else if (address_i == 8'd197) begin
      data_d[196:0] = data_q[196:0];
      data_d[197] = data_i;
      data_d[255:198] = data_q[255:198];
    end else if (address_i == 8'd198) begin
      data_d[197:0] = data_q[197:0];
      data_d[198] = data_i;
      data_d[255:199] = data_q[255:199];
    end else if (address_i == 8'd199) begin
      data_d[198:0] = data_q[198:0];
      data_d[199] = data_i;
      data_d[255:200] = data_q[255:200];
    end else if (address_i == 8'd200) begin
      data_d[199:0] = data_q[199:0];
      data_d[200] = data_i;
      data_d[255:201] = data_q[255:201];
    end else if (address_i == 8'd201) begin
      data_d[200:0] = data_q[200:0];
      data_d[201] = data_i;
      data_d[255:202] = data_q[255:202];
    end else if (address_i == 8'd202) begin
      data_d[201:0] = data_q[201:0];
      data_d[202] = data_i;
      data_d[255:203] = data_q[255:203];
    end else if (address_i == 8'd203) begin
      data_d[202:0] = data_q[202:0];
      data_d[203] = data_i;
      data_d[255:204] = data_q[255:204];
    end else if (address_i == 8'd204) begin
      data_d[203:0] = data_q[203:0];
      data_d[204] = data_i;
      data_d[255:205] = data_q[255:205];
    end else if (address_i == 8'd205) begin
      data_d[204:0] = data_q[204:0];
      data_d[205] = data_i;
      data_d[255:206] = data_q[255:206];
    end else if (address_i == 8'd206) begin
      data_d[205:0] = data_q[205:0];
      data_d[206] = data_i;
      data_d[255:207] = data_q[255:207];
    end else if (address_i == 8'd207) begin
      data_d[206:0] = data_q[206:0];
      data_d[207] = data_i;
      data_d[255:208] = data_q[255:208];
    end else if (address_i == 8'd208) begin
      data_d[207:0] = data_q[207:0];
      data_d[208] = data_i;
      data_d[255:209] = data_q[255:209];
    end else if (address_i == 8'd209) begin
      data_d[208:0] = data_q[208:0];
      data_d[209] = data_i;
      data_d[255:210] = data_q[255:210];
    end else if (address_i == 8'd210) begin
      data_d[209:0] = data_q[209:0];
      data_d[210] = data_i;
      data_d[255:211] = data_q[255:211];
    end else if (address_i == 8'd211) begin
      data_d[210:0] = data_q[210:0];
      data_d[211] = data_i;
      data_d[255:212] = data_q[255:212];
    end else if (address_i == 8'd212) begin
      data_d[211:0] = data_q[211:0];
      data_d[212] = data_i;
      data_d[255:213] = data_q[255:213];
    end else if (address_i == 8'd213) begin
      data_d[212:0] = data_q[212:0];
      data_d[213] = data_i;
      data_d[255:214] = data_q[255:214];
    end else if (address_i == 8'd214) begin
      data_d[213:0] = data_q[213:0];
      data_d[214] = data_i;
      data_d[255:215] = data_q[255:215];
    end else if (address_i == 8'd215) begin
      data_d[214:0] = data_q[214:0];
      data_d[215] = data_i;
      data_d[255:216] = data_q[255:216];
    end else if (address_i == 8'd216) begin
      data_d[215:0] = data_q[215:0];
      data_d[216] = data_i;
      data_d[255:217] = data_q[255:217];
    end else if (address_i == 8'd217) begin
      data_d[216:0] = data_q[216:0];
      data_d[217] = data_i;
      data_d[255:218] = data_q[255:218];
    end else if (address_i == 8'd218) begin
      data_d[217:0] = data_q[217:0];
      data_d[218] = data_i;
      data_d[255:219] = data_q[255:219];
    end else if (address_i == 8'd219) begin
      data_d[218:0] = data_q[218:0];
      data_d[219] = data_i;
      data_d[255:220] = data_q[255:220];
    end else if (address_i == 8'd220) begin
      data_d[219:0] = data_q[219:0];
      data_d[220] = data_i;
      data_d[255:221] = data_q[255:221];
    end else if (address_i == 8'd221) begin
      data_d[220:0] = data_q[220:0];
      data_d[221] = data_i;
      data_d[255:222] = data_q[255:222];
    end else if (address_i == 8'd222) begin
      data_d[221:0] = data_q[221:0];
      data_d[222] = data_i;
      data_d[255:223] = data_q[255:223];
    end else if (address_i == 8'd223) begin
      data_d[222:0] = data_q[222:0];
      data_d[223] = data_i;
      data_d[255:224] = data_q[255:224];
    end else if (address_i == 8'd224) begin
      data_d[223:0] = data_q[223:0];
      data_d[224] = data_i;
      data_d[255:225] = data_q[255:225];
    end else if (address_i == 8'd225) begin
      data_d[224:0] = data_q[224:0];
      data_d[225] = data_i;
      data_d[255:226] = data_q[255:226];
    end else if (address_i == 8'd226) begin
      data_d[225:0] = data_q[225:0];
      data_d[226] = data_i;
      data_d[255:227] = data_q[255:227];
    end else if (address_i == 8'd227) begin
      data_d[226:0] = data_q[226:0];
      data_d[227] = data_i;
      data_d[255:228] = data_q[255:228];
    end else if (address_i == 8'd228) begin
      data_d[227:0] = data_q[227:0];
      data_d[228] = data_i;
      data_d[255:229] = data_q[255:229];
    end else if (address_i == 8'd229) begin
      data_d[228:0] = data_q[228:0];
      data_d[229] = data_i;
      data_d[255:230] = data_q[255:230];
    end else if (address_i == 8'd230) begin
      data_d[229:0] = data_q[229:0];
      data_d[230] = data_i;
      data_d[255:231] = data_q[255:231];
    end else if (address_i == 8'd231) begin
      data_d[230:0] = data_q[230:0];
      data_d[231] = data_i;
      data_d[255:232] = data_q[255:232];
    end else if (address_i == 8'd232) begin
      data_d[231:0] = data_q[231:0];
      data_d[232] = data_i;
      data_d[255:233] = data_q[255:233];
    end else if (address_i == 8'd233) begin
      data_d[232:0] = data_q[232:0];
      data_d[233] = data_i;
      data_d[255:234] = data_q[255:234];
    end else if (address_i == 8'd234) begin
      data_d[233:0] = data_q[233:0];
      data_d[234] = data_i;
      data_d[255:235] = data_q[255:235];
    end else if (address_i == 8'd235) begin
      data_d[234:0] = data_q[234:0];
      data_d[235] = data_i;
      data_d[255:236] = data_q[255:236];
    end else if (address_i == 8'd236) begin
      data_d[235:0] = data_q[235:0];
      data_d[236] = data_i;
      data_d[255:237] = data_q[255:237];
    end else if (address_i == 8'd237) begin
      data_d[236:0] = data_q[236:0];
      data_d[237] = data_i;
      data_d[255:238] = data_q[255:238];
    end else if (address_i == 8'd238) begin
      data_d[237:0] = data_q[237:0];
      data_d[238] = data_i;
      data_d[255:239] = data_q[255:239];
    end else if (address_i == 8'd239) begin
      data_d[238:0] = data_q[238:0];
      data_d[239] = data_i;
      data_d[255:240] = data_q[255:240];
    end else if (address_i == 8'd240) begin
      data_d[239:0] = data_q[239:0];
      data_d[240] = data_i;
      data_d[255:241] = data_q[255:241];
    end else if (address_i == 8'd241) begin
      data_d[240:0] = data_q[240:0];
      data_d[241] = data_i;
      data_d[255:242] = data_q[255:242];
    end else if (address_i == 8'd242) begin
      data_d[241:0] = data_q[241:0];
      data_d[242] = data_i;
      data_d[255:243] = data_q[255:243];
    end else if (address_i == 8'd243) begin
      data_d[242:0] = data_q[242:0];
      data_d[243] = data_i;
      data_d[255:244] = data_q[255:244];
    end else if (address_i == 8'd244) begin
      data_d[243:0] = data_q[243:0];
      data_d[244] = data_i;
      data_d[255:245] = data_q[255:245];
    end else if (address_i == 8'd245) begin
      data_d[244:0] = data_q[244:0];
      data_d[245] = data_i;
      data_d[255:246] = data_q[255:246];
    end else if (address_i == 8'd246) begin
      data_d[245:0] = data_q[245:0];
      data_d[246] = data_i;
      data_d[255:247] = data_q[255:247];
    end else if (address_i == 8'd247) begin
      data_d[246:0] = data_q[246:0];
      data_d[247] = data_i;
      data_d[255:248] = data_q[255:248];
    end else if (address_i == 8'd248) begin
      data_d[247:0] = data_q[247:0];
      data_d[248] = data_i;
      data_d[255:249] = data_q[255:249];
    end else if (address_i == 8'd249) begin
      data_d[248:0] = data_q[248:0];
      data_d[249] = data_i;
      data_d[255:250] = data_q[255:250];
    end else if (address_i == 8'd250) begin
      data_d[249:0] = data_q[249:0];
      data_d[250] = data_i;
      data_d[255:251] = data_q[255:251];
    end else if (address_i == 8'd251) begin
      data_d[250:0] = data_q[250:0];
      data_d[251] = data_i;
      data_d[255:252] = data_q[255:252];
    end else if (address_i == 8'd252) begin
      data_d[251:0] = data_q[251:0];
      data_d[252] = data_i;
      data_d[255:253] = data_q[255:253];
    end else if (address_i == 8'd253) begin
      data_d[252:0] = data_q[252:0];
      data_d[253] = data_i;
      data_d[255:254] = data_q[255:254];
    end else if (address_i == 8'd254) begin
      data_d[253:0] = data_q[253:0];
      data_d[254] = data_i;
      data_d[255] = data_q[255];
    end else if (address_i == 8'd255) begin
      data_d[254:0] = data_q[254:0];
      data_d[255] = data_i;
    end
  end else begin
    data_d = data_q;
  end
end

always @(posedge clk_i) begin
  data_q <= data_d;
end

endmodule
